//dut
module dut(
  //...
  );
endmodule
